`ifndef PARAMETER_H_
`define PARAMETER_H_

// Parameter file

`define instruction_column 16 
`define data_column 16 
`define instruction_row 15
`define data_row 8 
`define filename "output.txt"
`define simulation_time #160

//this is to enable random input instruction
`define RANDOM_INSTRUCTION_INPUT

`endif
